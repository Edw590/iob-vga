assign im_pixel_x = pixel_x;
assign im_pixel_y = pixel_y;
assign rgb = im_rgb;
